LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY Deslocador IS 
 GENERIC(N: natural := 8);
 PORT(entrada	: IN  STD_LOGIC_VECTOR(N-1 DOWNTO 0);
		  saida		: OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0));
END ENTITY;

ARCHITECTURE comportamento OF Deslocador IS

FUNCTION desloca(ent : STD_LOGIC_VECTOR(N-1 DOWNTO 0)) RETURN STD_LOGIC_VECTOR IS
VARIABLE aux1 : STD_LOGIC_VECTOR(N-1 DOWNTO 0);
BEGIN
   aux1:=ent(N-3 downto 0)&"00";
	RETURN aux1;
END;

BEGIN
saida <= desloca(entrada);
END ARCHITECTURE;
